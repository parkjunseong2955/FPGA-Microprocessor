`timescale 1ns / 1ps

module tb_TOP();

// input
reg clk_ref; // reference clock
reg [3:0] sw; // switch 신호
reg [3:0] btn; // button 신호

//output
wire [1:0] seg_en; // SSD 활성화 신호
wire [6:0] seg_ab, seg_cd; // SSD 출력 신호
wire [3:0] led; //LED 출력 신호

always #4 clk_ref = ~clk_ref; // 125MHz clock 생성

// TOP module을 UUT로 호출 및 입출력 port 매핑
TOP uut(.clk_ref(clk_ref), .sw(sw), .btn(btn), .seg_en(seg_en), .seg_ab(seg_ab), .seg_cd(seg_cd), .led(led));

initial begin
    clk_ref = 0; btn = 4'b0000; sw = 4'b0000;  // initial value
#10              btn=4'b1000;                  // reset

// WRITE 동작 테스트
#10              btn = 4'b0001;                // S0 -> S1 (button[0]을 활성화)
#1000          btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                         sw = 4'b0001; // opcode: 1(wirte)
#10000         btn = 4'b0001;                // S1 -> S2
#5000          btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                       //sw = 4'b0000; // rd1: don't care
#10000         btn = 4'b0001;                // S2 -> S3
#5000          btn = 4'b0000;                // S3: 명령어 입력 3 (rd2)
#10000                         sw = 4'b0101; // rd2: 0101(5) 
#10000         btn = 4'b0001;                // S3 -> S4
#5000          btn = 4'b0000;                // S4: 명령어 입력 4 (wr)
#10000                         sw = 4'b0001; // wr: $1
#10000         btn = 4'b0001;                // S4 -> S5
#5000          btn = 4'b0000;                // S5: 실행
#10000         btn = 4'b0001;                // S5 -> S6
#5000          btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000         btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기 
#10000         btn = 4'b0000;                // button[1] 땜(다시 실행결과 2진수로 출력)
#5000          btn = 4'b1000;                // S6 -> S0 (idle 상태로 초기화)
#10000         btn = 4'b0000;                // S0

// ADD 동작(ADDI도 동일), ADDI에서는 rd2:I
#10              btn = 4'b0001;                // S0 -> S1
#1000          btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                         sw = 4'b1010; // opcode: 10(add)
#10000         btn = 4'b0001;                // S1 -> S2
#5000          btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                         sw = 4'b0001; // rd1: $1
#10000         btn = 4'b0001;                // S2 -> S3
#5000          btn = 4'b0000;                // S3: 명령어 입력 3 (rd2)
#10000                         sw = 4'b0010; // rd2: $2
#10000         btn = 4'b0001;                // S3 -> S4
#5000          btn = 4'b0000;                // S4: 명령어 입력 4 (wr)
#10000                         sw = 4'b0011; // wr: $3
#10000         btn = 4'b0001;                // S4 -> S5
#5000          btn = 4'b0000;                // S5: 실행
#10000         btn = 4'b0001;                // S5 -> S6
#5000          btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000         btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기 
#10000         btn = 4'b0000;                // butto[1] 땜(다시 실행결과 2진수로 출력)
#5000          btn = 4'b1000;                // S6 -> S0 (idle 상태로 초기화)
#10000         btn = 4'b0000;                // S0

// READ 동작
#10              btn = 4'b0001;                // S0 -> S1
#1000          btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                         sw = 4'b0010; // opcode: 2(read)
#10000         btn = 4'b0001;                // S1 -> S2
#5000          btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                         sw = 4'b0011; // rd1: $3
#10000         btn = 4'b0001;                // S2 -> S3
#5000          btn = 4'b0000;                // S3: 명령어 입력 3 (rd2)
#10000                       //sw = 4'b0100; // rd2: don't care 
#10000         btn = 4'b0001;                // S3 -> S4
#5000          btn = 4'b0000;                // S4: 명령어 입력 4 (wr)
#10000                       //sw = 4'b0001; // wr: don't care
#10000         btn = 4'b0001;                // S4 -> S5
#5000          btn = 4'b0000;                // S5: 실행
#10000         btn = 4'b0001;                // S5 -> S6
#5000          btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000         btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기 
#10000         btn = 4'b0000;                // button[1] 땜(다시 실행결과 2진수로 출력)
#5000          btn = 4'b1000;                // 상태 변환 S6 -> S0 (idle 상태로 초기화)
#10000         btn = 4'b0000;                // S0

// SUB 동작
#10              btn = 4'b0001;                // S0 -> S1
#1000            btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                          sw = 4'b1011;  // opcode: 11 (SUB)
#10000           btn = 4'b0001;                // S1 -> S2
#5000            btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                          sw = 4'b0001;  // rd1: $1
#10000           btn = 4'b0001;                // S2 -> S3
#5000            btn = 4'b0000;                // S3 : 명령어 입력 3 (rd2)
#10000                          sw = 4'b0010;  // rd2: $2
#10000           btn = 4'b0001;                // S3 -> S4
#5000            btn = 4'b0000;                // S4 : 명령어 입력 4 (wr)
#10000                          sw = 4'b0011;  // wr: $3
#10000           btn = 4'b0001;                // S4 -> S5
#5000            btn = 4'b0000;                // S5: 실행
#10000           btn = 4'b0001;                // S5 -> S6
#5000            btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000           btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기
#10000           btn = 4'b0000;                // button[1] 땜
#5000            btn = 4'b1000;                // S6 -> S0 (idle 상태로 초기화)
#10000           btn = 4'b0000;                // S0

// AND 동작
#10              btn = 4'b0001;                // S0 -> S1
#1000          btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                         sw = 4'b0101; // opcode: 5(and)
#10000         btn = 4'b0001;                // S1 -> S2
#5000          btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                         sw = 4'b0011; // rd1: $3
#10000         btn = 4'b0001;                // S2 -> S3
#5000          btn = 4'b0000;                // S3: 명령어 입력 3 (rd2)
#10000                         sw = 4'b0010; // rd2: $2 
#10000         btn = 4'b0001;                // S3 -> S4
#5000          btn = 4'b0000;                // S4: 명령어 입력 4 (wr)
#10000                         sw = 4'b0011; // wr: $3
#10000         btn = 4'b0001;                // S4 -> S5
#5000          btn = 4'b0000;                // S5: 실행
#10000         btn = 4'b0001;                // S5 -> S6
#5000          btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000         btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기 
#10000         btn = 4'b0000;                // button[1] 땜(다시 실행결과 2진수로 출력)
#5000          btn = 4'b1000;                // S6 -> S0 (idle 상태로 초기화)
#10000         btn = 4'b0000;                // S0

// SLL 동작
#10              btn = 4'b0001;                // S0 -> S1
#1000            btn = 4'b0000;                // S1 : 명령어 입력 1 (op)
#10000                          sw = 4'b1110;  // opcode: 14 (SLL)
#10000           btn = 4'b0001;                // S1 -> S2
#5000            btn = 4'b0000;                // S2 : 명령어 입력 2 (rd1)
#10000                          sw = 4'b0001;  // rd1: $1 (Shift할 값)
#10000           btn = 4'b0001;                // S2 -> S3
#5000            btn = 4'b0000;                // S3 : 명령어 입력 3 (rd2)
#10000                          sw = 4'b0011;  // rd2: Shift Amount (3)
#10000           btn = 4'b0001;                // S3 -> S4
#5000            btn = 4'b0000;                // S4 : 명령어 입력 4 (wr)
#10000                          sw = 4'b0010;  // wr: $2
#10000           btn = 4'b0001;                // S4 -> S5
#5000            btn = 4'b0000;                // S5: 실행
#10000           btn = 4'b0001;                // S5 -> S6
#5000            btn = 4'b0000;                // S6: done (실행결과 2진수로 출력)
#10000           btn = 4'b0010;                // button[1] 누르면 실행한 명령어 ssd에 표기
#10000           btn = 4'b0000;                // button[1] 땜
#5000            btn = 4'b1000;                // S6 -> S0 (idle 상태로 초기화) -> 상태만 초기화, 값은 그대로
#10000           btn = 4'b0000;                // S0
#100 $finish;
end

endmodule